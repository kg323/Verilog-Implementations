/*
Name: Kenneth Galindo
Class: ECE 526 Lab
Lab Report: #3
File Name: Lab3_1
*/

module dff (q, qbar, clock, data, clear);
	input clock, data, clear;
	output q, qbar;

	not #

endmodule
